module display_com(In,Out);
	input [3:0] In;
	output [13:0] Out;
	reg [13:0] Out;
	always @(*)
		case(In)
			4'b0000: Out=14'b11111111000000; //0
			4'b0001: Out=14'b11111111111001; //1
			4'b0010: Out=14'b11111110100100; //2
			4'b0011: Out=14'b11111110110000; //3
			4'b0100: Out=14'b11111110011001; //4
			4'b0101: Out=14'b11111110010010; //5
			4'b0110: Out=14'b11111110000010; //6
			4'b0111: Out=14'b11111111111000; //7  		   
			4'b1000: Out=14'b01111111111000; //8
			4'b1001: Out=14'b01111110011000;  //9
			4'b1010: Out=14'b01111110000010;  //10
			4'b1011: Out=14'b01111110010010;  //11
			4'b1100: Out=14'b01111110011001;  //12
			4'b1101: Out=14'b01111110110000;  //13
			4'b1110: Out=14'b01111110100100;  //14
			4'b1111: Out=14'b01111111111001;  //15

		endcase
endmodule
